package alu_pkg;

//standard UVM import & include

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "transaction_item.sv"
`include "alu_config.sv"
`include "alu_driver.sv"
`include "alu_sequence.sv"
`include "alu_sequencer.sv"
`include "alu_env.sv"
`include "alu_test.sv"

endpackage: alu_pkg
